interface test_if(
                    input logic clk, 
                    input logic rstn 
                    );
endinterface