`define WORD_SIZE 32
`define INST_SIZE 32

`define BYTE_SIZE 8
`define HALF_SIZE `WORD_SIZE/2

`define DM_DEPTH  256 //Data Memory depth
`define IM_DEPTH  256 //Instruction Memory depth

`define DM_FILE "mem.rv32i" //File tha initialize Data Memory
`define IM_FILE "Code_Examples/RV32I/I_Type_Test.rv32i" //File that initializes Instruction Memory

`define N_REG 32
//`define TEST