`timescale 1ns / 1ps
//`define TEST
//`define TEST_FILE//Test using the file functions
`define FPGA

module INSTRUCTION_MEMORY(
    output [31:0] o_Instruction,
    input [31:0] i_Addr
    );

	parameter HEIGHT = 76;//Memory height
	parameter FILE = "test2.r32i";

	reg [7:0] mem [HEIGHT-1:0];//Memory: Word: 1byte

	`ifdef TEST
	//This block is used for tests
	initial begin
		$readmemh(FILE, mem);//Initialize Memory
	end
	`endif

	`ifdef FPGA
	/*
		The instruction memory is initialized with the hexadecimal code generated by the assembler.
	It's used one C code (Mount.c) to generate this initilization.
	*/
	initial begin
		mem[0]='hE0;
		mem[1]='h06;
		mem[2]='hE0;
		mem[3]='h05;
		mem[4]='h00;
		mem[5]='h43;
		mem[6]='h00;
		mem[7]='h00;
		mem[8]='h08;
		mem[9]='h00;
		mem[10]='h00;
		mem[11]='h00;
		mem[12]='h08;
		mem[13]='h04;
		mem[14]='h00;
		mem[15]='h00;
		mem[16]='h1B;
		mem[17]='hF8;
		mem[18]='h1B;
		mem[19]='hFF;
		mem[20]='h37;
		mem[21]='hFF;
		mem[22]='h37;
		mem[23]='hFF;
		mem[24]='h37;
		mem[25]='hFF;
		mem[26]='h32;
		mem[27]='hFF;
		mem[28]='h68;
		mem[29]='hC1;
		mem[30]='h68;
		mem[31]='hC1;
		mem[32]='h60;
		mem[33]='h0A;
		mem[34]='h60;
		mem[35]='h0A;
		mem[36]='h68;
		mem[37]='h81;
		mem[38]='h68;
		mem[39]='h81;
		mem[40]='h68;
		mem[41]='h46;
		mem[42]='h68;
		mem[43]='h46;
		mem[44]='h1B;
		mem[45]='hFA;
		mem[46]='h32;
		mem[47]='h55;
		mem[48]='h60;
		mem[49]='h0A;
		mem[50]='h60;
		mem[51]='h0A;
		mem[52]='h47;
		mem[53]='hB0;
		mem[54]='h1B;
		mem[55]='hFA;
		mem[56]='h32;
		mem[57]='hAA;
		mem[58]='h60;
		mem[59]='h0A;
		mem[60]='h60;
		mem[61]='h0A;
		mem[62]='h47;
		mem[63]='hB0;
		mem[64]='hE7;
		mem[65]='hF4;
		mem[66]='h1B;
		mem[67]='hFD;
		mem[68]='h3D;
		mem[69]='h01;
		mem[70]='h1B;
		mem[71]='hED;
		mem[72]='hD7;
		mem[73]='hFD;
		mem[74]='h47;
		mem[75]='h70;
	end
	`endif

	assign o_Instruction = {mem[i_Addr+3], mem[i_Addr+2], mem[i_Addr+1], mem[i_Addr]};//One instruction has 32 bits


endmodule
