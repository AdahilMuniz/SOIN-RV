`define TESTE //Define for select test parts of code  
`define FPGA //Defines for select FPGA parts of code