//DEFINES
`include "../defines/ALU_CONTROL.vh"
`include "../defines/OPCODES_DEFINES.vh"
`include "../defines/PARAMETERS.vh"
`include "../defines/PROJECT_CONFIG.vh"

//RV32I Files
`include "ALU.v"
`include "ALU_CONTROL.v"
`include "DATA_MEMORY.v"
`include "DATAPATH.v"
`include "IMM_GENERATOR.v"
`include "INSTRUCTION_MEMORY.v"
`include "MAIN_CONTROL.v"
`include "REGISTER_FILE.v"
`include "DATAPATH.v"
`include "CORE.v"