/*************/
/***MACHINE***/
/*************/

/*Address*/
`define MISA_ADDR 'h301

/*Content*/
//MISA
`define MISA_MXL 2'h1
`define MISA_EXTENSION 26'h0000100