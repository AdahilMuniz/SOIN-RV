`define WORD_SIZE 32

`define DM_DEPTH  256 //Data Memory depth
`define IM_DEPTH  256 //Instruction Memory depth

`define DM_FILE "mem.rv32i" //File tha initialize Data Memory
`define IM_FILE "../../Code_Examples/RV32I/I_Type_Test.rv32i" //File tha initialize Instruction Memory

`define TEST