import types_pkg::*;

interface test_if(
                    input logic  clk, 
                    input logic  rstn,
                    input addr_t pc
                    );

endinterface